library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;  
-- Instruction Memory of the NYU-6463 Processor
entity Instruction_Memory is
port (
 pc: in std_logic_vector(31 downto 0);
 instruction: out  std_logic_vector(31 downto 0)
);
end Instruction_Memory;

architecture Behavioral of Instruction_Memory is
 type Instr_MEM is array (0 to 31) of std_logic_vector(31 downto 0);
 --R1=1,R2-=2.R3=3,R4=-2,R5=5
 constant instruction_data: Instr_MEM:=(
   -- AND: R1 and R2 -> R3  000000 00001 00010 00011 0 0000 010010 
   b"00000000001000100001100000010010", --pc=0
   -- ANDI: R1 and 3 -> R3  000011 00011 00001 0000000000000011 
   b"00001100011000010000000000000011", --pc=4
   -- OR: R1 or R2 -> R3  000000 00001 00010 00011 0 0000 010011 
   b"00000000001000100001100000010011", --pc=8
   -- NOR: R1 nor R2 -> R3  000000 00001 00010 00011 0 0000 010100
   b"00000000001000100001100000010100", --pc=12
   -- ORI: R1 or 3 -> R3  000100 00011 00001 0000000000000011 
   b"00010000011000010000000000000011", --pc=16
    -- Load word: MEM[R1+1] -> R3  000111 00011 00001 0000000000000001 (MEM[2] load to R3)
   b"00011100011000010000000000000001", --pc=20
    -- Store word: R1 -> MEM[R1+6]   101011 00001 00001 0000000000000110 (R1 store to MEM[3])
   b"10101100001000010000000000000110", --pc=24
   -- BLT: if R2 < R1, goto pc = PC+4+(1<<2)  001001 00001 00010 0000000000000001 (should not branch)
   b"00100100001000100000000000000001", --pc=28
   -- BEQ: if R2 = R1, goto pc = PC+4+(1<<2)  001010 00001 00010 0000000000000001 (should not branch)
   b"00101000001000100000000000000001", --pc=32
   -- BNE: if R2 != R1, goto pc = PC+4+(1<<2)  001011 00001 00010 0000000000000001 (should branch to pc = 40)
   b"00101100001000100000000000000001", --pc=36
   
   b"00000000000000000000000000000000", --pc=40
   -- JMP: goto pc = PC+4+(1<<2)  001100 00000 00000 0000000000000001 (should jump to pc = 52)
   b"00110000000000000000000000000001", --pc=44
   
   b"00000000000000000000000000000000", --pc=48
   -- ADD: R1 + R2 -> R3  000000 00001 00010 00011 0 0000 100000 (1+2=3)
   b"00000000001000100001100000100000", --pc=52
   -- ADDU: R1 + R4 -> R3  000000 00001 00100 00011 0 0000 100001 (1-2=-1)
   b"00000000001001000001100000100001", --pc=56
   -- ADDI: R1 + 5 -> R3  001000 00011 00001 0000000000000101 
   b"00100000011000010000000000000101", --pc=60
   -- DIVU: R5/R2 -> R30,R31 000000 00101 00010 11110 0 0000 011010  (5/2 =2...1) 
   b"00000000101000101111000000011010", --pc=64
   -- XRLR: R5 xor R2, lfrot 2 -> R3 000000 00101 00010 00011 0 0010 010000 ( (5 xor 2) <<2 ) 
   b"00000000101000100001100010010000", --pc=68
    -- RRXR: R5 rtrot 2, xor R2 -> R3 000000 00101 00010 00011 0 0010 010001 ( (5>>2 xor R2 ) 
   b"00000000101000100001100010010001", --pc=72
    -- LRAD: R5 lfrot 2 + R2 -> R3 000000 00101 00010 00011 0 0010 010101 ( (5<<2 + R2 ) 
   b"00000000101000100001100010010101", --pc=76
   -- SBRR: R5 - R2, rtrot 2 -> R3 000000 00101 00010 00011 0 0010 010110 ( (5-2, rr 2 )
   b"00000000101000100001100010010110", --pc=80
   
      -- DIVU: R5/R0 -> R30,R31 000000 00101 00000 11110 0 0000 011010  (5/0 =X...X) 
   b"00000000101000001111000000011010", --pc=84
   
   -- HAL: halt 111111 00000000000000000000000000
   b"11111100000000000000000000000000",--pc=88
   
   b"00000000000000000000000000000000",
   b"00000000000000000000000000000000",
   b"00000000000000000000000000000000",
   b"00000000000000000000000000000000",
   b"00000000000000000000000000000000",
   b"00000000000000000000000000000000",
   b"00000000000000000000000000000000",
   b"00000000000000000000000000000000",
   b"00000000000000000000000000000000"
  );
begin
 instruction <= instruction_data(to_integer(unsigned(pc(31 downto 2))));

end Behavioral;